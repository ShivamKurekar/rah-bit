/* encode the mipi frame to send to processor */
module rah_encoder (
    input                                   clk,
    input                                   vid_gen_clk,

    input [TOTAL_APPS-1:0]                  send_data,
    input [TOTAL_APPS-1:0]                  wr_clk,
    input [(TOTAL_APPS*DATA_WIDTH)-1:0]     wr_data,

    output [TOTAL_APPS-1:0]                 wr_fifo_full,
    output [TOTAL_APPS-1:0]                 wr_almost_fifo_full,
    output [TOTAL_APPS-1:0]                 wr_prog_fifo_full,

    output reg                              mipi_rst = 1,
    output                                  mipi_valid,
    output [DATA_WIDTH-1:0]                 mipi_data,
    output                                  hsync_patgen,
    output                                  vsync_patgen
);

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="ipecrypt"
`pragma protect encrypt_agent_info="IP Encrypter LLC, http://ipencrypter.com, Version: 23.7.0"
`pragma protect author="Vicharak"
`pragma protect author_info="Vicharak Computers Pvt Ltd"

`pragma protect key_keyowner="Efinix Inc."
`pragma protect key_keyname="EFX_K01"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_block
jpy8GXfSwqVrA+hZP2vzpqPNiboqZT0nmvFEz+hcO4PJMht1g696FuMUV4FWkLT5
1ismz1ODTFxQOot8gEmBhSVjwwHzEwjWw2g4bxYWahsPinOaIouX1x/Yw979t/5b
MfO+KhztEbLsCji8dz+i72/lesUhpSgQiuQk54GKxXG3msm4wjRgPRRs8HxtxsXY
QbaTQ3mrvxoHyanj0YLG9yOA8wisDNMlf5GNpYsfyiHoV98evWEb/9d47e0xxsOF
7UyTrQ7XoVSifO7RpqaD4sFXhkrDtu3GbQ+b2RIGfoeGNS1iiE3yfqmaAIKsBCGe
zd1aSEFCyno+O5z38811Rg==

`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_block
jOp53wT121w7MNjyeL6Nk1hOs3YWv84UXlgzFhhyxcgMFk5IUkQvqQwyv0rl9Wvp
2rUe90mPwZMeQ8eV/BphiCSfaRfx7swQGCRL5H8erp3IoTpcSlrc1WnG6NATfk3U
dssGT28eZy+Uf5lnSE2cpaNlQUtjF92I0VuotQaVE3Q=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=9890)
`pragma protect data_block
uXJ4CfwWzmEOYICH5Erman+J0vFVlJpPW15d4rQQj7odUJJcx3t+g4NXvsHjYVIZ
bOSDJbVnWRRjjdSqCi33iV6x8sMQyjPrV4WRKzUbrlaMAx8HTPgAymsf9D5h0BfR
nZP/DamqmPkVeZnIMxv1n/++bcVU61FXIEB10Z4rcm9DZp5jZVx44smgiup1fKe0
LbTTAlBp+MQP71tlUQar/9r1DGqzBdmOVeuxH6FgeXt61Jlyzrj0TZKZ9Z1XXyyN
jEjcwbLWleTJZ/F66UUf9HXYIK9sYoVvnI4QFMY1fSU2iQyZiPqB7vuq1FF+wk8j
bjQKIR4BCfLEucdd65QeeEzvx8Tsx2nepGUaz/YGYng/LKkgCybv+UYCzkBZZCCT
kdNyu84WfmJlra3ZuP2osPS9KeJwSICVvg/Y+Z5FkE+HhISMR13ek42dL4nKN6zr
qacyWEStkgj+rfCnIpP/mEaAIGNmkkzL2y3zHKHZ0JyNGyfkLC7YNGX6aI5a6uUl
j3oo5Byfjb/cG2TeMk0K7gJxhpGL9P8kvtoHJ+c6y/gn0lXPhbMZS4TALTlaPDC8
cROIjl44YgO5rAgwc2cc0r+hAN++UDEexe3mpp4Vzk8nVvaU6SMRf2BghS5A888u
kVNuyKc4YDdevHZ8EFOfPo/vxtRodLzkccnQhEcStQ6xsLUJbEoZJg42zd7hu1R4
as08dDxBOKvuikyEKrCvw7NJCUISTwVjlv98fjqrXNlFNYelvsqhZ2VxYRDNBp25
LlnTviKQAdGJub5BV7QOZJ2F4hdG0F8btBdR3nL3Kn9gF9X1zQtxnOSFkKIGBlmg
7asqsI0Eik23Bkv77S7I3S0BgIPe4KFzKeBtZqRb0zbSTa/Gl+pwg1QopzNByrfG
bDy6+cUjTDN4Nh+iIuxRXPSqNMzBV7aj8OkM3WZ6cn7nltCcXP7ObZ5m7gNyKKxV
1dOJZegbAJ6GGqb1Mg6ZoLKIgNkYuTlYJl6jf5tsrRb0hhxJver0LwcBP02ECv4A
FjMaZHwZt9aE7E4PiHmCtouNKBMedeA3uFPBSF0LGbcD8SJNvopDS/zBLcMdGWqh
faiTz4FBxvXHIk7feX5q9oe/LTxaq1NwnO3vaBbmX/yAVfizBV767bpv6q9hpGCj
pTqtbw44+tIiSVTP4rKNhd719vZKB4P802TKU55Ag0kzHl7CXwo388IrtO6JFfIe
LIq8cRxfr5BPmp3adfaPHH2lV8RyKRVYnWUZJbncbjuO3mpio/MNGtKwLIF25Tu+
0m0UITQR4ZEGdOZIcrov9goCDkYRXYGf4zY4jjljTO6wlsecAnUyWFuevq1yfIAb
IRLZBbxev9c/smbKDeKv+UGhYhHLtdE43EPju/mRKSEf3S1s3RG02m1uGf8JMpMs
qNpJ8wXPpkRvYJ7HX3jQLf3huLnLGBCIbVDcowPX+vZdi/Pe24RPjhFrq9ZoHrIm
eCuFJ+WQbGuGFkERLNTZRG0DNjxMoIOITtBZPNK10SWKRsod9dR2OwjvD65Xhkuq
bslf5Vuppuc3BTrf++RhyXEjMr6f4kUyMx3XtGSYfYCbzKc46bRi3baU5JLsOF0g
LF34dIS75kQ5J8Wli5hhQ2Qlgp2j7hfQfGsvlQdEoAbYeJYuxwCwa5B8T+ml1M9U
WP4LEAI3FLnilwHmrbfmH6uM4LU0QiI5yZB3RdFZOc38kZUNNX3vZE/FHvxXdXZd
PhzzAVV29m/k53MxzC8X36BnyHCVJG+S1dZqgWPyG08fGpA++D3wMaqvG4W+mxFm
9GvcPMA/4xZnjBMWVzrEQzw5BGFpv6aYszrfbWri+L6RLO7bSj8JtgDSNsjwK6nb
md/3zJD6FdOdcbIS8l4eTl8G2OrvPSnMcVYjgJVYYaCDvjBLVnyNvhMzSD7kaW29
JEZ7vbJjb53/gc5S0nQB/PgmWOC90/3mTvODFCxfGT10dB3IlPZ/zaMyt46bw71Y
SX9AtK/aQI3Si/B3hAF9fzCjISoFTMCZnA64wNuTois7w5S8U9ROJ/dKJLvuJMMw
2DJYz6VscvcNrN79VbnzHxwANhP9Ai1WeacUGVSPBH14VBJ+evFihTqaeOe3bLze
pt29OBfs2VmTVTdN7m6i8J/FAgK2rHCfSCqzrG731InhgBaqVd9GslAtFx32FzMW
/iGroi6e1VP6YceHHmTVioQGuwjG/m0VnzDuTQY6FpwqvSBTZlUbG6B+/9q3inzQ
a6D3B3J6fHlS1mgyVUc9jllhyR23X/iya6+ugVRHtSwEs/6nmxQv5vZCQ4Yvt0UN
xQ7DQTna90k0Z+42bWKbQw57M85hkr7Vc9XzlyXVNaBF4fJpjg2uGe2qT2a8HVgn
V33ynIXUo1xZ7ZxKcnmkguTQOTyjlF7ip7CqWz5UAFFcSxATB51eC53PXvOwl1kd
jTlSyNAYv30pdmb/LbJlYLmYA2UFDBzk6VVwcqRErOzX/cepczCXkE43m4t0JRe3
oh6nUzqJ02FnoqA0cVGnmEp3k3ZhPVvLzUwWBkDdFj+ZwRo2FsEhEvXfI/LdrT5C
COHuKN1RkbzVx+UKQUEbkMEScwdGpz2yvfyY0OGgu456mR18h4KtImHObJMzOToq
29+TLopn1/DgW8orbBuFOzIcqdoIY+pCHATM48lkd8K5PplKNCMVUzYwgxCyDruL
9W5tKhMG4nb+MgmZptICCwDPlMpfrEVu2tkAoBpxbMua8Q2KN2E0bQ2QpRA3SwUC
MjV7k4VlyTfF3DQOr1ja44cCvaXWoBUUkNR8d1UyrPWktanTkeopZY7iP2SrAYoW
JjlK7M7wAjPNE6tdEvNUZqHtBgJCsKO2pMyn78IOk8P2ZImKo9M0vw/KtOvEKrja
xn4qsGE/VSmqx6bkuq/1FPqJs9RBZPf+mbrrE9Gnfh5zjzmihKlF7Ry5eZ2WwkcF
ZptKl44PsdvYRaYZKuFA5KMbjWRZ0aiwJqs8tP6nRkceMdbFoKjs6LeYwBV69W8x
3kSj0ukFz79tcQyy+2sOigbWYJ8uy69GsHDJgNpavBTpnvNtI4fAsSCYELzgLMV2
xn1ledGoQmm2gwvltgLRHSyWKKhDwT70n0dfD1fhGEkqsMZnmXIXrjv16Ivc2O80
MPxhOwpQzmZoARMu5fAE4uSroWLS6PcGY9xaRu+Bz1h3LOMeUIRd7osEbzto1gq8
iDKf/hYIITkHTFdr/Gn7YLFLgczSzzpepliyQSQsW0xAiQP8Qd+3K+2kfM8wMGun
4nl0HEcuj86RHGqO1LhFbsr/hxt4iVSeDoxAc9g3qFxz5M99zlIskjgb2nagVeJD
5+Su2pinJEdR4LtFZsEXAID1Ds1Mlgi3LPjyqZsO+Fvt0wWWGlzU3n1WNszfoF0w
lUdK5XfC/J+7E92med2YFZByatA0YS3pHem0pzkKXsN4qYiMQQjtztVT0tkpCjx+
Bk1jLL3eh5WGwiVqwJr6oa7PXV4rNtzt1FX6R+UO8d7iYtLxztYAnA/eJ+kFUw/E
vcePfX11eoI4t3ogtphW8hPgwA0Tba1B7Ff55m36voiRAz6MnceLGEHA6lhHtXZ7
E/CFC8ElfJSCfEDCfx+w0Y8cItxZpwvpTCZROJaqS6MHiyHY1a48/vkw6RrbhDFt
tEpj9EcfmVtmg2HtqTMdHZuaT2cm6Nr89288cCKozzq85NyhmpCUnko5M4A2r107
uLgi+DKDzRIjhaIFWxBF4HxR3cj6t0KuxpkPLt1whbAm5FZdE22SyoNKd/pGDGx1
ZdBRyfD+86PRkMV8pW28x0OMqymxfxwjwOKA90we0BEaxhDD37CFm8QbwE08vCTU
8luZHcXYIJQgPT+yXZH9lrCdlwgNqVoXSewQlAgZW3XJK9EipoFrz/lZEsU1vB8Z
cVdXO49Nc7XC5BSlow7RuvR2RC3uPkzhsvNBqOq9JITUnS10Bmi7BlMTozlzCokL
wwGTd6t/emmfTmbXukX3OzUwT6QKtbr9mwpnb7LdTWT+1e9DG9dmA7uv9dZxxoTM
JPClmJBj+0aXbv6lhXka6WnSnRmhBgImEEot/okYbS0SCSsLUc8GwJt89cgoZ25v
Ai0nJSWtVT3twutpUIbiIIpEeRpKsUhEYOznmrtkcDW88a+obccqnH8tcE3tr0by
V7Z/1wdcqrJMpS4VLEr6eal72DpwiFinsZleEHSR+T22kZ7RVGHBcKhowBVje9Zz
jWMJeiV2DNf3XNj+im6FlCFnNVdpGY/tTo6JJn4S5rahtRqXQpLJzh0f6zqSoZRC
FmyCi+u+PBkP0eE1RkuSiaemEVHYw7slGzqRRTPCeFUalaTPYx7kJAY+zE62fhXj
Mejtqq6GMh/WpQq/VZV5V/e3iwgV4SxyDzNzwcI97IGFfuou3iHylcJZVakYM/TI
Ha4q3HdfogqUugw/kY9Q6VjyHDTjbbpwODnyzS/1bzbH0Dsp9fexQ7I8Z1IntloS
qr2rFF3h3a4tDXR+CEYaS7Vlg7ubiRK75+wE7RN+FszxwHOYxWobJS9ATs1ZlnKi
CIkrW2P6KiE5yhCsJcOFJlqVdigA52qPeLyYNW06iAd4oeTq1uUHP69DJqYRhY0m
A4RzjK+pcAmOzVIPVD/nZeTvqOl5PponvC9cesTvgyFb9KhhG+ts9xaPkNZwguIm
KkpF4qCUMFWIgae3tQeDa12m4UFHMX5nZxEMdTGH2tRd2QauTnKsfng+VGS3b4lf
yhgPg4ooliDFxZZ9FqNvHxIXL+beCvPs3V2/7l7EuhDdZgjNGgILZbsFeUrqxEMA
S4aJHKSxyd8FcQOciE0SKLiZ5pwKlD4K6KP2Le/hqrSAAOBnhpfDyK+Rx1alZNct
yddQnsfyeaUKOwm+2osbS6cl5VTnnSv3/J4QxZRTbN+hiPm6OKGxTKKkb9YQvKba
e1AAI/b2OTNV8DVv8ON7flTYqb0Gut8sV8AusrKsvqvQ8fBk06CMHMN0Qk2euI3F
lwAqmQJRTFJBtpFcudHKC7tE51fv8ommzcYR4GKMQY4P9pA8gr5U1Ymn1MSKvyTd
MM58VXGffFAjdT9fIL8uAx8L4+ay2Dhl8WAAkTbpG6BQvgfz66U/GlQoIHLzxy1J
KmoSNBd7liGAs/N+YqDTZrMt5O/UXZhFKPx3djTgoGi/Wg/2wOQrMBrsc05gbl7p
nkoiIj0+Gmg24H5Qrz/BHNJnjGOcht+MPL6+o5oIeFUznXWu/d3ECiu5FFs+POM2
c4ej6pBsFVeyp04ZbyHf8xgzGdpxuwqnmIFI1T94858EXFSW7GdAFvW7lYgnzBOv
iJnRyyJkxgz0BqcW2KDaHcQfoPqPEOkB6KyUJGX+7sq9FoSRREyzP0KBrOSsr4PY
UF+RQ5CjGGvGQbc9KacCbx07E8y38WxQ8ODryWrWvR3g+CobNB6bSuYBAIwOuJPi
WDcBhjnez4x1s/dPzU7YxaygNdlgNWDQbc5T3hvxzYGaXxxpVtPTJ6fU+sGWObon
cQJJueJqX5Jwqk+KW1kEG46pELVqmYUBrB/uiPtBy1mGcBuQgDBme2I0S8RDAacR
GJFREmx3Zk6xLg8AgfT3UK99pO02pA8T0VraHPN0E2+zwvk4MMrqnIWjvMQ3wBPz
YcoVnhtsFxUjD8Uz+kKL+XYvcWzEomoG5Wh1Uqy48EzmmJiox4RzdTC6z45GwiDy
K3JdHG3deVxL9OZL9GCcayIW+7vqE6uBZ9ZYZYOV81vBgPinRwR25IjBvG1oKtHd
iG0zXIDyj01P5Zm8QmxEhdCxfw5hVFAq+RyWnhg86iSvvDuQ2yD7V1X7YqCehsqX
9OZkxiaW/gp+ua/uKCp2ukXekh4Bx8yT6GGTtRqc+jLA9WMJwJ5a/acUKklnrmBy
Xk37xHaNU68hhZdOUZY3e/fHM3d+wZ+Q5H+b666WHZq8Zlb4YyHY2FXhxZ6MROOs
aDAkyP6UaoHuBjzoMpS0dt3ny12gtIy4GE/2KBJDbROZLF6YCNNFhw0FJ4pCZALd
RcTSZCP+st7FUJZoBQ8xBJ3CYGLe9KEWbppO5iEa1ebf/2R7fdNHwBU2iVA3kGZx
bvKiQ9WnxKoQSeYBMGhglbkVZcdPs+8bm12H8fAKkRiaryDuc6QT3I0GBnXWA40U
5B+4srdrZzWEbSbHOS/qDtWPwKOTx10AFvDLk3+JYHw/c7UTNT01xj5XaE0z0ddn
g8tlCTM7sHhr8QwFe1VthiKS+iH7DA+ANS8dd7fpYB5PuKY74avdzAZi8iXHnfBB
UMZyBeVRVMmtqYoC7IpOI1NZ6a/nKs0zqy4XCQLvsPbNmz70y0TW19JrXuOq/sm6
EBe27ZwFS9fUPYiF4xD1qe5Jqq7pZVji2SmzNBnf6HnieZUoxoUqOUaRMZuOoI6B
nvh0b8dUSqo2n5aPqjJNBreEhiZys8U9aAotxYlZB/MqHZJUWTc9NHaTwhPGqvXH
VM8bzzTbY4MQ6U6plyNSCvsti79uG7qYMigEhsYW9m6eR0Das+vOlxurUBboYrYz
1U/nCtBF5T/louKvt4hPZw+ZEMedC+HR2AKp3gNi8vPR53QBCJCDHKAVOZrZfu+2
cWyOSRCJaqvinCceTJPW2ngdyKtLfnyTQQa8EkrSkAL8cdU7O8ul1PCws/uAFiIx
h3YyIZnk+a5eRj/hTWL1V9+u9Rhf1lU6pv1ufoowgHKOG5Kl5SA8KRVpPCvAiv5i
kXzQGMBzg5c4+9KDlbSCdyQSmypvqn9RiY5cAKx6ySEo2sr8+TvE8FWbWINBKZnR
9JS6b+7Tqbezw+NgYTSeEC2FI5FiLLoXy4yM5e6SgYKRDTz9ko95PtaMtw6XHlg3
zhWabGx/p7v/tAx1SjgWHjqlpfhW8W6q33ews9wGTDTobwSZgt8rNYAL5KUUzUjJ
MNJGdaxaPde21JovBtmWAAoYIQjQGd43bqmoUSHN4RhW/dxCZDjT6ctSbobISM6S
7i2bD5fNILxCW/E8cORo6BJ5/txO2A4n4mY0hTnISu0SlVdcElT49aC7Xb2K/7CC
C9MeWE843cI6OG9Ni6aC87rPQSxwj25YsLGQoVhd5FpALGEyCmSqd3sWFBGUP8B0
GM4L84g36Uo2qlsf2aEg6Iw3AW/p98zf7aPnLxeRwl1qhI7hUasxiW1XRdAFEM/9
QtIPZA4bgKnMe9OsNacabnJZr0lJM/sU7IlZi0DGAbYx7zFPiwHlOLtYmMrmean1
A3Y8YPc58OQ053GjukX+m7bHP9mLlqxDDzGpEhPkBrebpqrXW/NXYDDkLJ8ISTbs
wEbPPxwY0TUd5yVCfSGsLorgtT7rNyqTaDyLOSHKtf0zuKVxD2aG+pMGEc5hDBmF
r1mC5Oj1PoXl3SsC3fQ1MGpPhVTKL7Jut/9r7B1tP8oJaMbERe5TCWyJcb943ojL
C9jtZOlzTv3TL7ixVL6lcy/ZBGmK/buuGHUwDyW4HYk9qlMaDXfx1CE+9WAQPlRW
A+Jl70pAySGHorwcxH80Xo4G1/J2aWwE5oK+QMTwMTEESZAPN+jW5cwZrLjAvOGO
KamVw85tOTXt2Y34b0Kw/JVlvyd4xTliBHo5XAp/oVW+uf6bLB+CRDU7IpWJsg+S
EH7pmbZh3uiiyESAAkJuChLgRC5E5/8O/hN3kFZ0fH6mV41Pg36sSE6Pa0tSsD3R
qoF5DokusErKOC20aGaoXDFquxP9yjxkkCy3QwqrPj428Y1ukcMjF+0z82CVMz6U
8FNYRz/8I5BRhqRAgul4N3kyz6qiuyZEnGoq3qYMf9/zgLbS0jcgwGIl02QiS77R
pBKBOMIiUlvtDXK6u0nYX6+6xBocBG/HZBE6/ennNsJpktjHZ/hIjZNQBRS3NCz/
qjav1yVgowUHM62yz5sFHpOH3iYDwmz44NQHBuIVq1KjgKYcNptECpMeIiBCGmaY
8Ls2F3l9m52kdvkirj1X+Gd8yJZHIN0QkkprX7bcpRO2VngVgVJhJe5U3pPOPgO8
issPgRRzuwY4I7yMDODt0mGjmLj8ydLTea4hudoll7onCp+k0LTgGIxGxQLdY1XX
vwQJ/WvHnkRyEQWstbIrvB4nYAP8tdJr2augJMTyhOri5m3bltNgI4pZhZjBQbft
KlJn3mt0JZaWGIWdPrmUiGDKFDfG0EiifRRXqHk5fHyXVkvBdKgjiwX4THAOwvBA
B3KywZxce0ttb6OIIabox27zrnfkfOa5TXRvnBP57egv5DyhnQk8nXAjDoNkYmyK
11BgAsxPh0oFWXuCzSRT7VMDdqWLlG+W7msTbi00i2a0Phd/NuLIh++wJLrlnkgm
ziTkhAYHuIP5PFi12TQM7zHKaOJx6WjJ0JiKOXcyQlMZKZad3QVBGNFMYjEm/fBw
qqjodwfVCtZ0lz8n+I1RQdcdfJThB8eYJGB8HHPizzlR1IqCq3xKjxWu6L3LN+e2
c/29KigqVoYqncJob0BRX62IbipqEy4qQGnJpXV8CNkjD/3Blnf4aMsH3rXCRco2
bDb50uD9nRsT+r06hBkczXHpRbMwTtxilI+GTgPJWpHHiKwN2ISYqlp6ujhzKzKt
BL4e/indAfi3ZVOcxdQJcpKHsAUl5argA2+j/mqSMSZj98y+OHLNQ2lTJufCxIE0
1iP2Yi1nDRmdpCRM4mt1/4ZQmaLm9jA52RR7MZpybziQWSAvTsnW92qKiKCtFFC1
7p6P6YSRgOHFCMrAm/F3JbcPU1ZAkfoYgDSvRXFG6fnMqnxucZ7ap7HFdcNWf1rs
mRO2msaylNOC8Do6b+WimlKpz3FV/+r97SP1Wd9S7eVnX0pHHhkIHnYTqd9wOEef
D4Vb2VoGqzG7KM1cx0SDXWp8U6hIl4hLzxHE3UUeiBtI0WrLRaw5esf+wcDhNYbN
tk7yzae22TFDCaMIrFHS+A+Wtd9UV27bQBvT+T+kQOJOURT0UjdZUPnab3pcJJry
YwJYTTE8caA+37jPEj/uNPaBkNYDFfZWPcffpNEtZCfz5mhGw/TiFqZfXZ0Zk9tp
/+1zGoQD04Mbq4+4zlzT9m+aNr6XTlZpC9AexVKxGdHEfNx4yg2wXCRZe96m8TFF
WgIkquZutDcKdwycMhqv6cS9KfU1aXURbie7TZ5hR49ro6I4hmfJt0AR9+uUMjcZ
bFnbe9ZBS7lE4FdOKCvSpdPpYkMAIyHw579HyinIvQuPv86JaqBufZ2d7b55PWZ0
y0fpKEnBv4X/cyRiejom8Cx4jMgYh2em7yP2Jtvn9HfgHjHYkMnu0i7ld+ZxCyK4
xFa2fw4h0Sq3aYtU43Ann9kfAA3RDRM73NknS7yu+YC7C5pN2eEKgpb+TGzKSnEa
vbPrr53Pi+CBS9ItEvnSQOr+/wL2j93eu0TA/S20r6wey2IcRbX/a8TFQijOd7Z9
2BGE57zxh3HgKu/sbH0V9zPd5AAo3btVwBeZ9IVawMDLg2VjjPS4N2zCNrG68hyn
jTbsPX830R/SfOv8H4iQPJZWaDXJuU06TRpwzgkbzV1XM0B0nhRr/Jny1YJXiDd1
pOiYTYtpLJZJav9/UhIKVL0ISJvS//yALnxGcWmd9ZHqQp9s1LQGRFEUqitUxhgR
gpbB4Lk50sbs9lD8oOt6sC69dwlPKhjpSdA1qGfF77RWaGSbqvRFeW/2H+DuqyOI
ajcqCmfKdEFLILiF2oEXeO6MoC+XpbecNz3wB4JKrnrqNM3p5ec6TrvrMK8+h6qX
aNffHMJ354lxbfEcwtja5FtmIr94qHk3pfAdE7Qv+cITr0YWwqbrkWdnPaqDgsYg
rmXwszBPH8hEN6Rg1MWkHJJuGDIg6urPgtDjOKABEZvqBrqVVyxRtgnLj7NGqvkP
LVqthj6D5pcyAhyIFvdmi1ihnNHgXLfp4sz8uWhIpc3BPX4U9nEPQ5KX538NszXT
NUPS9b9nL05fkwmHL4TG+EUPgimbPig4et/5gbELIM3vfabB7Wzt/XXYHMy8sbhd
bCtlxgU0CueuvenjoGU8iRdToh3Xcwc+UseZVLCm35bdGJOTQ6zRqHrTyVdzTiVX
a3tDwMna5Rs7X6i1DAUfiQF3DyJgdX7S5jRAv2cnkMFdmzcFY2FOMxHA8E0i0wQY
g6n5vKd0vIkW97i7vYBLIjxzaFZLvzCO6QjTjOc6vDVeW1R6sFVGoemVEn2igGGw
aE8ANqpLdIdnaDZVPOeoN9Az8D/7bm4QldSnVCMx1ZE2G2TjRiaZmv0P1XgiIerx
SsShaSNzF4zHnb+R6PY+xqwUoKstwRwAS07uP41q3U8LqNWZDYyCYZoo69IGH0lR
3VUsUx3kxzf73d5zUz/KekUKHTcSCEZuIKroCxergDiuVG90VbCLe9mTCLWdWqvI
iQQM9oJrfHiVfQrtb5sdf6IGzur8h6XwjJQI7tCWsM9ajFA9RgRGYP4v/lKouF6K
xVRl3jD7UpGmgRoxYR7+QLStZ3hCvV8qELN98TNhsw+56Bc+pkYb1tDGCvvWznk7
8Q4boJPpb6/CzSnJlxyk60PqNFOvQrc/hjhndv2ERETQGTTgYQtuSGggavU467am
uGnRuyfTDdTyD6YtQqxaWBeEAhLQo8UQQltUI38JJIaBu4k0l5ooRIxSpY2rS90c
j63geKKhrsMlIkhBi5aGEP6YAMfN8rRBh2bY6MMRLP4Ocfd2p7jh5xC7IT7Chckp
GPbKbffrq4bau6BW6CRXGFJQX+Jbh2Hjj5NLjsybg+Xk+C1kA+kkZhjUnv1gjSI8
hO4Ex5xZI0aTJEbmZXsPGdg7tfWq5auqL5mLEXj+x83vyXgNtDtZCi8QE7z1M/0z
i8VJK0NG5FZguDd+PJRv+7Zam42gUJicErpsmzrC6ThJgAu1XC2N9XImpOhk1pJT
ZQhq5GeubPQ8DWNvhVVDiuFoxwrrkvLUj678zIXXHBF6bPdOQzljTUexuxGiLeEm
mWVna0r5/aFXYNFdisZI1w8sGFCAE4YZibY419Fr9wQnVM35xuG9WYpUiN3iB9i9
icckuZMg544dzl3Qsr72t5QSk1BHu1t/esKfeqF7elNKDX4Y5LTr+xB05y+LnRrR
u8udLhfTWwZcbs6jtRtU+Fdb2lZLGPvtlO8+/HM5SfMJnmr+o9NLKFkQe/wKM6xc
Kp38TyiOzKfX4+JIbO2uxPWtxZ48GLaJ0pDuEYIuKinkPySVo1XCdJ4UVIJUhQBF
ksFcXr9oeNShBytmLiRZ3iLXbhFe9OqMNlfZtO1Roz9hI4jp23ZNRKAAXatoITkx
C7WIWpJJ0/NVcYb9sISelWiICmlIXYXTSMnuLTiIUN1l0rVjHo2BOgD/nyrIAqTI
G+rxHqhHmhxolb9RwL389AfqZkh9tfjJLtLGIA6Lnmu73gjfVRU63LGBQB6hTJnT
J31JC40YhGbutlxxfSSt92bxBxbzcq9E4uFwzeAgpFR14YuallZxjDmbJfw/eUhL
sb1Zn5MCX3gFLa0BE/Pj6NVuhYizmzuVnkeD3U/S6/U7vPKq+qJM9f7nLxUc0tz0
Hcx5FPsQGvgUbey8xm1MBUEJpnw7hfJvn1nLHM5brcWtnGf4GjP2ryA6gkFDFVfx
1VQWTn+YgyXNmQrFZTrsIojL/zyjCVmyGyE32TIaWabj2gs7VQZyS4cg1iYiyNzx
zLjU75PUrZ/3q+ChrYS+kNcuvy4/ePwDHZ0K2kAuTlb4vWlm6yZytscieG4g47yb
qSYp/76lB3LXyjD/dzz0UogOvr3g4bAkeUsNyDYPjZlvRTCxQhi4mF/NX1dOQmZu
0DBq0ZHpJqytubVsUEfKDY1aWjaIjAs+sEqdawypWwfBVAQj/yNQ1lPMTB7WxphF
Ri/bf+sX5wz2oEpgQbyspvRhjKHrnO1ubeyjJmq6Qqh/9BP0LKfIK176FDrtt47q
WQD+07IjFc/nT1wLIGfSKZoWgP1qoS3k6FLmkal8q2WWkiqFuZXbVAnMlzHIF/+q
aejg8X+26SI/iJwxizEXv2uPqyrTwXXVRv6uC70x1il87m6lxkxctu9L+zsd52Xq
ACAcm0XPrguxs9z52Y8URJ0//gdntcMkATBObyVf6sRKoR0aMtV5Ddtkfhe771m3
Il0I/VcftwwVElpgKc9enNvgoWSMSPHQadlI/no9wMu2LzCYXrgza4EDnbm6QY9S
CzU03F6VBRMVOvW9G/zBuRh0SrobRgdXzw3mPsa1NPj8Eay++XfcE9rla/GZKklx
uX592RKL3j/rgMNgxX8gtS1jSzEl668fESV8xfZAKLxs2Ocpx3Y3ob8EYszzwi4o
HargPyObrAjIkQaus1iWbHahvMs9GrizwTu70/njbkv8Dlf3YVCVk9vrDCduIlv1
5b33M6gmrxmP2Y+NLpSVasFrZs58fXn0Zwk91ZKg02uPLSe+fPUI8IQCWC+mJK+n
XHsuzOQFi67F1YUjJJxMo/AXiXrAawq0uTJ0sd7tZbs0AOUP/qBOTtOJCL5nUV65
Dwk+uv+2o0l6neP1733vtFQtxIBBMAdc0eLO9/RKqevMrLCj5pI3pBrOjuR8Ruwu
+wApN7e90Hz4pLNa8AjuXdyFbzn51uNnQWk2ArHlWqVCb4kU1oLPvetHmoMks7O3
7SHrQDzv4omIpgUq0G7fBdSf7xNA6o5uF87GE886S4yhzhBdbF472Q3q6DrPUOyD
LI8YC9QqGRczAcpRuIZP4vJCntJOK3FAUCKR6OPkMDRq/Sx5atjrSGs+gmMA0Gd+
GB/Ir2iP/SKzEdcSTk24clEo5QiiOCtwcc3KzEWIpjXIakUyYLBHFJMTM6RM8UxA
RQ6cx6v8Wj8I0HRLrY/KVMFLMsUrXcS9axAXnCBQ9xeSqGLOserNdgNZkY5v1UJM
Mx8Q6lWRHouSMJOMHPxFUQJ6rPb8MLwqqMGnXNoyqtd0wQuPC8dBS6BFankR5i3O
qEOT5DpDcpf1OvXQvRyiTxl69L3+Ermz0x6Ab55VNMfKZraOPQlcysYJ47mPwGPr
aqYWGLr0ySDOLB2EEApuUrjeS4nltTY5SVnuZlfy9RXeNr2DcWkfAGonh/vgQlsi
IGON4SGrHaNU/KyogBHTtKQ35joa73VwGucbAvwg8f3N/HK6xBvKOdNiEoJDMKBh
fkf8JesSOO/JgrOpxSxdGF4M5aN4OHADfFW4FNaNpS6UPUW/KC9TtGagP1UMeibQ
J19tMMKlKiVubs8HMserBA==
`pragma protect end_protected

endmodule
